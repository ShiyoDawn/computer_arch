library verilog;
use verilog.vl_types.all;
entity fadd_vlg_vec_tst is
end fadd_vlg_vec_tst;
