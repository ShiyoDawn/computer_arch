library verilog;
use verilog.vl_types.all;
entity alucomb_vlg_vec_tst is
end alucomb_vlg_vec_tst;
