library verilog;
use verilog.vl_types.all;
entity hadd8_vlg_vec_tst is
end hadd8_vlg_vec_tst;
