library verilog;
use verilog.vl_types.all;
entity alusys_vlg_vec_tst is
end alusys_vlg_vec_tst;
