library verilog;
use verilog.vl_types.all;
entity dec3_8_vlg_vec_tst is
end dec3_8_vlg_vec_tst;
