library verilog;
use verilog.vl_types.all;
entity dec2_4_vlg_vec_tst is
end dec2_4_vlg_vec_tst;
