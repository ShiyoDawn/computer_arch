library verilog;
use verilog.vl_types.all;
entity alu_ROM_vlg_vec_tst is
end alu_ROM_vlg_vec_tst;
