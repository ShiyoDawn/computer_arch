library verilog;
use verilog.vl_types.all;
entity sh1c_vlg_vec_tst is
end sh1c_vlg_vec_tst;
