library verilog;
use verilog.vl_types.all;
entity ALU8_181_vlg_vec_tst is
end ALU8_181_vlg_vec_tst;
