library verilog;
use verilog.vl_types.all;
entity selector_vlg_vec_tst is
end selector_vlg_vec_tst;
