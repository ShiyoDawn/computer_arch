library verilog;
use verilog.vl_types.all;
entity addsub8_vlg_vec_tst is
end addsub8_vlg_vec_tst;
