library verilog;
use verilog.vl_types.all;
entity add8_vlg_vec_tst is
end add8_vlg_vec_tst;
