library verilog;
use verilog.vl_types.all;
entity regg_vlg_vec_tst is
end regg_vlg_vec_tst;
