library verilog;
use verilog.vl_types.all;
entity addsub8 is
    port(
        Co              : out    vl_logic;
        Ci              : in     vl_logic;
        M               : in     vl_logic;
        A               : in     vl_logic_vector(7 downto 0);
        B               : in     vl_logic_vector(7 downto 0);
        S               : out    vl_logic_vector(7 downto 0)
    );
end addsub8;
