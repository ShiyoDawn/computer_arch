library verilog;
use verilog.vl_types.all;
entity ks_test_vlg_vec_tst is
end ks_test_vlg_vec_tst;
