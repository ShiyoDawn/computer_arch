library verilog;
use verilog.vl_types.all;
entity sel2g_vlg_vec_tst is
end sel2g_vlg_vec_tst;
