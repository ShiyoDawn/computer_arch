library verilog;
use verilog.vl_types.all;
entity sel4g_vlg_vec_tst is
end sel4g_vlg_vec_tst;
