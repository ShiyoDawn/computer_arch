library verilog;
use verilog.vl_types.all;
entity ramsub_vlg_vec_tst is
end ramsub_vlg_vec_tst;
