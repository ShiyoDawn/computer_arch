library verilog;
use verilog.vl_types.all;
entity hadd_vlg_vec_tst is
end hadd_vlg_vec_tst;
